`define FEATURE_ICACHE_STAT
// Width of byte enable for a given data width
`define EVAL_BE_WIDTH(DATAWIDTH) (DATAWIDTH/8)


`define NB_CORES  8
`define SH_NB_CACHE_BANKS  2
